library ieee;
use ieee.std_logic_1164.all;

entity execute is
end entity;

architecture execute_arq of execute is


begin
end architecture;